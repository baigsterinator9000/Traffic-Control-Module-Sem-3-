NET "Clock" LOC = "p1"|IOSTANDARD=LVCMOS33; # CMOD-P35 - GCK2, Global Clock Input

#System level constraints
Net Clock TNM_NET = Clock;
Timespec TS_Clock = PERIOD Clock 10us; #adjust to suit Clock, 10us->100kHz

#Reset pin
NET "Reset" LOC = "p30"|IOSTANDARD=LVCMOS33; # CMOD-P18 - GCK2, Global Set/Reset
Net "Reset" TIG;

NET "CarEW" LOC = "p33"|IOSTANDARD=LVCMOS33; # CMOD-P24 - GTS0, Global Tristate Control
NET "CarNS" LOC = "p34"|IOSTANDARD=LVCMOS33; # CMOD-P25 - GTS1, Global Tristate Control

NET "PedEW" LOC = "p36"|IOSTANDARD=LVCMOS33; # CMOD-P26 - I/O
NET "PedNS" LOC = "p37"|IOSTANDARD=LVCMOS33; # CMOD-P27 - I/O

NET "LightsEW<1>" LOC = "p39"|IOSTANDARD=LVCMOS33; # CMOD-P29 - I/O
NET "LightsEW<0>" LOC = "p40"|IOSTANDARD=LVCMOS33; # CMOD-P30 - I/O

NET "LightsNS<1>" LOC = "p41"|IOSTANDARD=LVCMOS33; # CMOD-P31 - I/O
NET "LightsNS<0>" LOC = "p42"|IOSTANDARD=LVCMOS33; # CMOD-P32 - I/O

NET "LEDs<0>" LOC = "p18"|IOSTANDARD=LVCMOS33; # CMOD-P9 - I/O
NET "LEDs<1>" LOC = "p19"|IOSTANDARD=LVCMOS33; # CMOD-P10 - I/O
NET "LEDs<2>" LOC = "p20"|IOSTANDARD=LVCMOS33; # CMOD-P11 - I/O
NET "LEDs<3>" LOC = "p21"|IOSTANDARD=LVCMOS33; # CMOD-P12 - I/O
NET "LEDs<4>" LOC = "p22"|IOSTANDARD=LVCMOS33; # CMOD-P13 - I/O
NET "LEDs<5>" LOC = "p23"|IOSTANDARD=LVCMOS33; # CMOD-P14 - I/O
NET "LEDs<6>" LOC = "p27"|IOSTANDARD=LVCMOS33; # CMOD-P15 - I/O
NET "LEDs<7>" LOC = "p28"|IOSTANDARD=LVCMOS33; # CMOD-P16 - I/O